module mac_tb;
endmodule
